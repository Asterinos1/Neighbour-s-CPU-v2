library IEEE;
use IEEE.STD_LOGIC_1164.all;

package arr_vector5 is
	type arr_v5 is ARRAY(NATURAL RANGE<>) OF STD_LOGIC_VECTOR(4 downto 0);
end package arr_vector5;