library IEEE;
use IEEE.STD_LOGIC_1164.all;

package matrices is
	type MATRIX is array(natural range<>) of std_logic_vector(31 downto 0);
end matrices;